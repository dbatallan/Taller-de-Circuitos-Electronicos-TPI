** Profile: "SCHEMATIC1-RegulacionDeCarga"  [ C:\Users\Lionheart\Documents\GitHub\Taller-de-Circuitos-Electronicos-TPI\Checkpoint 1\Version 2.5 - Limitador de Corriente Basico  - Etapa de ganancia de tencion intermedia\Orcad\Version 2-5-PSpiceFiles\SCHEMATIC1\RegulacionDeCarga.sim ] 

** Creating circuit file "RegulacionDeCarga.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Lionheart\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC DEC PARAM RVAL 0.0001 1k 30 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
